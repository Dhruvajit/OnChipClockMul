PLL CIRCUIT
V2 Fclkin 0 PULSE(0 1.8 10p 10p 10p 100n 200n)
V4 VIN 0 1.8
XX9 Fclkin output DOWN UP pfd_cmos_baker_nand_not
XX4 DOWN UP vco_input chargepumpf
C1 vco_input 0 146p
C2 vco_input N001 500p
R1 N001 0 500
XX5 0 VIN vco_input vco_out vco_f
XX1 vco_out VIN N003 frequencydividerby2new
XX2 N003 VIN N002 frequencydividerby2new
XX3 N002 VIN output frequencydividerby2new



*BLOCK SYMBOL DEFINITION
*--------------------------------------------------
*PHASE FREQUENCY DETECTOR
.subckt pfd_cmos_baker_nand_not Frequency_in Frequency_VCO down up
XX1 vdd Frequency_in 0 N005 not
XX2 vdd N002 0 N003 not
XX3 vdd N003 0 N004 not
XX4 vdd N001 0 up not
XX5 vdd Frequency_VCO 0 N012 not
XX6 vdd N009 0 N014 not
XX7 vdd N014 0 N015 not
XX8 vdd N013 0 down not
XX9 N001 N005 vdd 0 N002 nand_2input
XX10 N002 N007 vdd 0 N006 nand_2input
XX11 N006 N008 vdd 0 N007 nand_2input
XX12 N008 N010 vdd 0 N011 nand_2input
XX13 N011 N009 vdd 0 N010 nand_2input
XX14 N012 N013 vdd 0 N009 nand_2input
XX15 N004 N006 N008 0 vdd N001 nand
XX16 N008 N010 N015 0 vdd N013 nand
XX17 N008 vdd 0 N006 N002 N009 N010 nand_4input
V1 vdd 0 1.8
.include osu018.lib
.ends pfd_cmos_baker_nand_not

*-------------------------------------
*FREQUENCY DIVIDER BY 2
.subckt frequencydividerby2new clock vdd Q
M1 Q_bar clock_bar N002 0 nfet l=.18u w=.18u
M2 N002 clock Q_bar vdd pfet l=.18u w=.54u
M3 N004 N002 0 0 nfet l=.18u w=.18u
M4 vdd N002 N004 vdd pfet l=.18u w=.54u
M5 N002 clock N003 0 nfet l=.18u w=.18u
M6 N003 clock_bar N002 vdd pfet l=.18u w=.54u
M7 N003 N004 0 0 nfet l=.18u w=.18u
M8 vdd N004 N003 vdd pfet l=.18u w=.54u
M9 N004 clock N001 0 nfet l=.18u w=.18u
M10 N001 clock_bar N004 vdd pfet l=.18u w=.54u
M11 N001 clock_bar Q_bar 0 nfet l=.18u w=.18u
M12 Q_bar clock N001 vdd pfet l=.18u w=.54u
M13 Q N001 0 0 nfet l=.18u w=.18u
M14 vdd N001 Q vdd pfet l=.18u w=.54u
M15 Q_bar Q 0 0 nfet l=.18u w=.18u
M16 vdd Q Q_bar vdd pfet l=.18u w=.54u
M17 clock_bar clock 0 0 nfet l=.18u w=.18u
M18 vdd clock clock_bar vdd pfet l=.18u w=.54u
.include osu018.lib
.ends frequencydividerby2new

*-------------------------------------
*CHARGE PUMP
.subckt chargepumpf DOWN UP CP
M1 N003 UP 0 0 nfet l=.18u w=.18u
M3 N005 DOWN 0 0 nfet l=.18u w=.18u
M4 VDD DOWN N005 VDD pfet l=.18u w=.54u
M5 VDD UP N003 VDD pfet l=.18u w=.54u
M7 N003 0 N001 N001 nfet l=.18u w=.18u
M8 N006 VDD N005 N006 pfet l=.18u w=.54u
M9 N005 0 N006 N006 nfet l=.18u w=.18u
M10 N004 N006 N004 N004 nfet l=.18u w=.18u
M11 0 VDD VDD 0 nfet l=.18u w=.18u
M12 N004 DOWN 0 0 nfet l=.18u w=15u
M13 CP VDD N004 N004 nfet l=.18u w=.18u
M14 N001 VDD N003 N001 pfet l=.18u w=.54u
M15 N002 UP N002 N002 pfet l=.18u w=.54u
M16 VDD N001 N002 VDD pfet l=.18u w=45u
M17 N002 0 CP N002 pfet l=.18u w=.54u
M18 0 0 VDD VDD pfet l=.18u w=.54u
V1 VDD 0 1.8
.include osu018.lib
.ends chargepumpf

*-------------------------------------
*VOLTAGE CONTROL OSCILLATOR
.subckt vco_f GND VDD Vin_vco Osc
M7 Vp Vn GND 0 nfet l=.18u w=.18u
M8 Vp Vp VDD VDD pfet l=.18u w=.90u
XU1 osc_fb N001 Vp Vn VDD 0 cs_inv
XU2 N001 N002 Vp Vn VDD 0 cs_inv
XU3 N002 N003 Vp Vn VDD 0 cs_inv
XU4 N003 N004 Vp Vn VDD 0 cs_inv
XU5 N004 N005 Vp Vn VDD 0 cs_inv
XU6 N005 next Vp Vn VDD 0 cs_inv
XU19 next osc_fb Vp Vn VDD 0 cs_inv
XU22 osc_fb Osc inv_20_10
R2 Vn Vin_vco 1
.include osu018.lib
.ends vco_f

*-------------------------------------
*PFD - 2 INPUT NAND
.subckt not vdd vin ground out
M1 vdd vin out vdd pfet l=.18u w=.36u
M2 out vin ground ground nfet l=.18u w=.18u
.include osu018.lib
.ends not

*-------------------------------------
*PFD - 2 INPUT NAND
.subckt nand_2input va vb vdd ground out
M1 out va N001 ground nfet l=.18u w=.36u
M2 N001 vb ground ground nfet l=.18u w=.36u
M3 vdd va out vdd pfet l=.18u w=.36u
M4 vdd vb out vdd pfet l=0.18u w=.36u
.include osu018.lib
.ends nand_2input

*-------------------------------------
*PFD - 3 INPUT NAND
.subckt nand va vb vc ground vdd out
M1 out va N001 ground nfet l=.18u w=.54u
M2 N001 vb N002 ground nfet l=.18u w=.54u
M3 N002 vc ground ground nfet l=.18u w=.54u
M4 vdd va out vdd pfet l=.18u w=.36u
M5 vdd vb out vdd pfet l=.18u w=.36u
M6 vdd vc out vdd pfet l=.18u w=.36u
.include osu018.lib
.ends nand

*-------------------------------------
*PFD - 4 INPUT NAND
.subckt nand_4input out vdd ground va vb vc vd
M1 vdd va out vdd pfet l=.18u w=.36u
M2 vdd vb out vdd pfet l=.18u w=.36u
M3 vdd vc out vdd pfet l=.18u w=.36u
M4 vdd vd out vdd pfet l=.18u w=.36u
M5 out va N001 ground nfet l=.18u w=.72u
M6 N001 vb N002 ground nfet l=.18u w=.72u
M7 N002 vc N003 ground nfet l=.18u w=.72u
M8 N003 vd ground ground nfet l=.18u w=.72u
.include osu018.lib
.ends nand_4input

*-------------------------------------
*STAGES IN VCO
.subckt cs_inv In Out Vp Vn VDD GND
M1 N002 Vn GND 0 nfet l=.18u w=.18u
M4 N001 Vp VDD VDD pfet l=.18u w=.54u
M3 Out In N001 VDD pfet l=.18u w=.54u
M2 Out In N002 0 nfet l=.18u w=.18u
C1 Out 0 1f
.include osu018.lib
.ends cs_inv

*-------------------------------------
*INVERTER OF VCO
.subckt inv_20_10 In Out
M1 Out In 0 0 nfet l=.18u w=.18u
M2 N001 In Out N001 pfet l=.18u w=.54u
V1 N001 0 1.8
.include osu018.lib
.ends inv_20_10

*-------------------------------------

*Model Statements
.include osu018.lib
.model NMOS nfet
.model PMOS pfet


.tran 1ns 10u

*Control Statements
.control
run
plot V(Fclkin)+10 V(output)+8 V(UP)+6 V(DOWN)+4 V(vco_input)+2 V(vco_out)

.endc
.end

