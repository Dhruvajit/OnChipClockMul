title
V2 Fclkin 0 PULSE(0 1.8 10p 10p 10p 100n 200n)
V4 VIN 0 1.8
XX9 Fclkin output DOWN UP pfd_cmos_baker_nand_not
XX4 DOWN UP vco_input chargepumpf
C1 vco_input 0 146p
C2 vco_input N001 500p
R1 N001 0 500
XX5 0 VIN vco_input vco_out vco_f
XX1 vco_out VIN N003 frequencydividerby2new
XX2 N003 VIN N002 frequencydividerby2new
XX3 N002 VIN output frequencydividerby2new



*BLOCK SYMBOL DEFINITION
*--------------------------------------------------
*PHASE FREQUENCY DETECTOR
.subckt pfd_cmos_baker_nand_not Frequency_in Frequency_VCO down up
XX1 vdd Frequency_in 0 N005 not
XX2 vdd N002 0 N003 not
XX3 vdd N003 0 N004 not
XX4 vdd N001 0 up not
XX5 vdd Frequency_VCO 0 N012 not
XX6 vdd N009 0 N014 not
XX7 vdd N014 0 N015 not
XX8 vdd N013 0 down not
XX9 N001 N005 vdd 0 N002 nand_2input
XX10 N002 N007 vdd 0 N006 nand_2input
XX11 N006 N008 vdd 0 N007 nand_2input
XX12 N008 N010 vdd 0 N011 nand_2input
XX13 N011 N009 vdd 0 N010 nand_2input
XX14 N012 N013 vdd 0 N009 nand_2input
XX15 N004 N006 N008 0 vdd N001 nand
XX16 N008 N010 N015 0 vdd N013 nand
XX17 N008 vdd 0 N006 N002 N009 N010 nand_4input
V1 vdd 0 1.8
.include osu018.lib
.ends pfd_cmos_baker_nand_not

*-------------------------------------
*FREQUENCY DIVIDER BY 2
.subckt frequencydividerby2new clock vdd Q
M1 Q_bar clock_bar N002 0 nfet l=.18u w=.18u
M2 N002 clock Q_bar vdd pfet l=.18u w=.54u
M3 N004 N002 0 0 nfet l=.18u w=.18u
M4 vdd N002 N004 vdd pfet l=.18u w=.54u
M5 N002 clock N003 0 nfet l=.18u w=.18u
M6 N003 clock_bar N002 vdd pfet l=.18u w=.54u
M7 N003 N004 0 0 nfet l=.18u w=.18u
M8 vdd N004 N003 vdd pfet l=.18u w=.54u
M9 N004 clock N001 0 nfet l=.18u w=.18u
M10 N001 clock_bar N004 vdd pfet l=.18u w=.54u
M11 N001 clock_bar Q_bar 0 nfet l=.18u w=.18u
M12 Q_bar clock N001 vdd pfet l=.18u w=.54u
M13 Q N001 0 0 nfet l=.18u w=.18u
M14 vdd N001 Q vdd pfet l=.18u w=.54u
M15 Q_bar Q 0 0 nfet l=.18u w=.18u
M16 vdd Q Q_bar vdd pfet l=.18u w=.54u
M17 clock_bar clock 0 0 nfet l=.18u w=.18u
M18 vdd clock clock_bar vdd pfet l=.18u w=.54u
.include osu018.lib
.ends frequencydividerby2new

*-------------------------------------
*CHARGE PUMP
.subckt chargepumpf DOWN UP CP
M1 N003 UP 0 0 nfet l=.18u w=.18u
M3 N005 DOWN 0 0 nfet l=.18u w=.18u
M4 VDD DOWN N005 VDD pfet l=.18u w=.54u
M5 VDD UP N003 VDD pfet l=.18u w=.54u
M7 N003 0 N001 N001 nfet l=.18u w=.18u
M8 N006 VDD N005 N006 pfet l=.18u w=.54u
M9 N005 0 N006 N006 nfet l=.18u w=.18u
M10 N004 N006 N004 N004 nfet l=.18u w=.18u
M11 0 VDD VDD 0 nfet l=.18u w=.18u
M12 N004 DOWN 0 0 nfet l=.18u w=15u
M13 CP VDD N004 N004 nfet l=.18u w=.18u
M14 N001 VDD N003 N001 pfet l=.18u w=.54u
M15 N002 UP N002 N002 pfet l=.18u w=.54u
M16 VDD N001 N002 VDD pfet l=.18u w=45u
M17 N002 0 CP N002 pfet l=.18u w=.54u
M18 0 0 VDD VDD pfet l=.18u w=.54u
V1 VDD 0 1.8
.include osu018.lib
.ends chargepumpf

*-------------------------------------
*VOLTAGE CONTROL OSCILLATOR
.subckt vco_f GND VDD Vin_vco Osc
M7 Vp Vn GND 0 nfet l=.18u w=.18u
M8 Vp Vp VDD VDD pfet l=.18u w=.90u
XU1 osc_fb N001 Vp Vn VDD 0 cs_inv
XU2 N001 N002 Vp Vn VDD 0 cs_inv
XU3 N002 N003 Vp Vn VDD 0 cs_inv
XU4 N003 N004 Vp Vn VDD 0 cs_inv
XU5 N004 N005 Vp Vn VDD 0 cs_inv
XU6 N005 next Vp Vn VDD 0 cs_inv
XU19 next osc_fb Vp Vn VDD 0 cs_inv
XU22 osc_fb Osc inv_20_10
R2 Vn Vin_vco 1
.include osu018.lib
.ends vco_f

*-------------------------------------
*PFD - 2 INPUT NAND
.subckt not vdd vin ground out
M1 vdd vin out vdd pfet l=.18u w=.36u
M2 out vin ground ground nfet l=.18u w=.18u
.include osu018.lib
.ends not

*-------------------------------------
*PFD - 2 INPUT NAND
.subckt nand_2input va vb vdd ground out
M1 out va N001 ground nfet l=.18u w=.36u
M2 N001 vb ground ground nfet l=.18u w=.36u
M3 vdd va out vdd pfet l=.18u w=.36u
M4 vdd vb out vdd pfet l=0.18u w=.36u
.include osu018.lib
.ends nand_2input

*-------------------------------------
*PFD - 3 INPUT NAND
.subckt nand va vb vc ground vdd out
M1 out va N001 ground nfet l=.18u w=.54u
M2 N001 vb N002 ground nfet l=.18u w=.54u
M3 N002 vc ground ground nfet l=.18u w=.54u
M4 vdd va out vdd pfet l=.18u w=.36u
M5 vdd vb out vdd pfet l=.18u w=.36u
M6 vdd vc out vdd pfet l=.18u w=.36u
.include osu018.lib
.ends nand

*-------------------------------------
*PFD - 4 INPUT NAND
.subckt nand_4input out vdd ground va vb vc vd
M1 vdd va out vdd pfet l=.18u w=.36u
M2 vdd vb out vdd pfet l=.18u w=.36u
M3 vdd vc out vdd pfet l=.18u w=.36u
M4 vdd vd out vdd pfet l=.18u w=.36u
M5 out va N001 ground nfet l=.18u w=.72u
M6 N001 vb N002 ground nfet l=.18u w=.72u
M7 N002 vc N003 ground nfet l=.18u w=.72u
M8 N003 vd ground ground nfet l=.18u w=.72u
.include osu018.lib
.ends nand_4input

*-------------------------------------
*STAGES IN VCO
.subckt cs_inv In Out Vp Vn VDD GND
M1 N002 Vn GND 0 nfet l=.18u w=.18u
M4 N001 Vp VDD VDD pfet l=.18u w=.54u
M3 Out In N001 VDD pfet l=.18u w=.54u
M2 Out In N002 0 nfet l=.18u w=.18u
C1 Out 0 1f
.include osu018.lib
.ends cs_inv

*-------------------------------------
*INVERTER OF VCO
.subckt inv_20_10 In Out
M1 Out In 0 0 nfet l=.18u w=.18u
M2 N001 In Out N001 pfet l=.18u w=.54u
V1 N001 0 1.8
.include osu018.lib
.ends inv_20_10

*-------------------------------------
*Model Statements

.model nfet NMOS (LEVEL=8 VERSION=3.2 TNOM=27 TOX=4.1E-9 XJ=1E-7 NCH=2.3549E17 VTH0=0.3823463 K1=0.5810697

+            K2=4.774618E-3 K3=0.0431669 K3B=1.1498346 W0=1E-7 NLX=1.910552E-7 DVT0W=0 DVT1W=0 DVT2W=0

+            DVT0=1.2894824 DVT1=0.3622063 DVT2=0.0713729 U0=280.633249 UA=-1.208537E-9 UB=2.158625E-18

+            UC=5.342807E-11 VSAT=9.366802E4 A0=1.7593146 AGS=0.3939741 B0=-6.413949E-9 B1=-1E-7 KETA=-5.180424E-4

+            A1=0 A2=1 RDSW=105.5517558 PRWG=0.5 PRWB=-0.1998871 WR=1 WINT=7.904732E-10 LINT=1.571424E-8 XL=0

+            XW=-1E-8 DWG=1.297221E-9 DWB=1.479041E-9 VOFF=-0.0955434 NFACTOR=2.4358891 CIT=0 CDSC=2.4E-4 CDSCD=0

+            CDSCB=0 ETA0=3.104851E-3 ETAB=-2.512384E-5 DSUB=0.0167075 PCLM=0.8073191 PDIBLC1=0.1666161 PDIBLC2=3.112892E-3

+            PDIBLCB=-0.1 DROUT=0.7875618 PSCBE1=8E10 PSCBE2=9.213635E-10 PVAG=3.85243E-3 DELTA=0.01 RSH=6.7 MOBMOD=1

+            PRT=0 UTE=-1.5 KT1=-0.11 KT1L=0 KT2=0.022 UA1=4.31E-9 UB1=-7.61E-18 UC1=-5.6E-11 AT=3.3E4 WL=0 WLN=1

+            WW=0 WWN=1 WWL=0 LL=0 LLN=1 LW=0 LWN=1 LWL=0 CAPMOD=2 XPART=0.5 CGDO=7.08E-10 CGSO=7.08E-10 CGBO=1E-12

+            CJ=9.68858E-4 PB=0.8 MJ=0.3864502 CJSW=2.512138E-10 PBSW=0.809286 MJSW=0.1060414 CJSWG=3.3E-10 PBSWG=0.809286

+            MJSWG=0.1060414 CF=0 PVTH0=-1.192722E-3 PRDSW=-5 PK2=6.450505E-5 WKETA=-4.27294E-4 LKETA=-0.0104078

+            PU0=6.3268729 PUA=2.226552E-11 PUB=0 PVSAT=969.1480157 PETA0=1E-4 PKETA=-1.049509E-3)


.model pfet PMOS (LEVEL=8 VERSION=3.2 TNOM=27 TOX=4.1E-9 XJ=1E-7 NCH=4.1589E17 VTH0=-0.3938813 K1=0.5479015

+            K2=0.0360586 K3=0.0993095 K3B=5.7086622 W0=1E-6 NLX=1.313191E-7 DVT0W=0 DVT1W=0 DVT2W=0 DVT0=0.4911363

+            DVT1=0.2227356 DVT2=0.1 U0=115.6852975 UA=1.505832E-9 UB=1E-21 UC=-1E-10 VSAT=1.329694E5 A0=1.7590478

+            AGS=0.3641621 B0=3.427126E-7 B1=1.062928E-6 KETA=0.0134667 A1=0.6859506 A2=0.3506788 RDSW=168.5705677

+            PRWG=0.5 PRWB=-0.4987371 WR=1 WINT=0 LINT=3.028832E-8 XL=0 XW=-1E-8 DWG=-2.349633E-8 DWB=-7.152486E-9

+            VOFF=-0.0994037 NFACTOR=1.9424315 CIT=0 CDSC=2.4E-4 CDSCD=0 CDSCB=0 ETA0=0.0608072 ETAB=-0.0426148

+            DSUB=0.7343015 PCLM=3.2579974 PDIBLC1=7.229527E-6 PDIBLC2=0.025389 PDIBLCB=-1E-3 DROUT=0 PSCBE1=1.454878E10

+            PSCBE2=4.202027E-9 PVAG=15 DELTA=0.01 RSH=7.8 MOBMOD=1 PRT=0 UTE=-1.5 KT1=-0.11 KT1L=0 KT2=0.022 UA1=4.31E-9

+            UB1=-7.61E-18 UC1=-5.6E-11 AT=3.3E4 WL=0 WLN=1 WW=0 WWN=1 WWL=0 LL=0 LLN=1 LW=0 LWN=1 LWL=0 CAPMOD=2 XPART=0.5

+            CGDO=6.32E-10 CGSO=6.32E-10 CGBO=1E-12 CJ=1.172138E-3 PB=0.8421173 MJ=0.4109788 CJSW=2.242609E-10 PBSW=0.8

+            MJSW=0.3752089 CJSWG=4.22E-10 PBSWG=0.8 MJSWG=0.3752089 CF=0 PVTH0=1.888482E-3 PRDSW=11.5315407 PK2=1.559399E-3

+            WKETA=0.0319301 LKETA=2.955547E-3 PU0=-1.1105313 PUA=-4.62102E-11 PUB=1E-21 PVSAT=50 PETA0=1E-4 PKETA=-4.346368E-3)

.tran 1ns 5u

*Control Statements
.control
run
plot V(vco_input)

.endc
.end

